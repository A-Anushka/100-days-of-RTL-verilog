module uni_ga(output y,input a,input b);
nand(y,a,b);
endmodule
