module d_to_bcd_tb( );
reg [9:0] y;
wire [3:0] a;
d_to_bcd a1 (a,y);
initial
begin
 #0  y=10'b0000000000;
 #50  y=10'b0000000001;
 #50  y=10'b0000000010;
 #50  y=10'b0000000100; 
 #50  y=10'b0000001000;
 #50  y=10'b0000010000;
 #50  y=10'b0000100000;
 #50  y=10'b0001000000; 
 #50  y=10'b0010000000;
 #50  y=10'b0100000000;
 #50 y=10'b1000000000;
#50 $finish;
end
endmodule
