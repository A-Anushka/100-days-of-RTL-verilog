module mux_4to1_tb( );
reg i0,i1,i2,i3;
reg s0,s1;
wire y;
mux_4to1 a1 (y,s0,s1,i0,i1,i2,i3);
initial 
begin
#0 s1=0;s0=0;i0=1;i1=0;i2=0;i3=0;           //s1 s0 = 0 0 --> y= i0
#50 i0=0;i1=1;i2=0;i3=0;                        
#50 i0=0;i1=0;i2=1;i3=0;
#50 i0=0;i1=0;i2=0;i3=1;

#50 s0=1;i0=1;i1=0;i2=0;i3=0;               //s1 s0 = 0 1 --> y= i1
#50 i0=0;i1=1;i2=0;i3=0;
#50 i0=0;i1=0;i2=1;i3=0;
#50 i0=0;i1=0;i2=0;i3=1;

#50 s1=1;s0=0;i0=1;i1=0;i2=0;i3=0;          //s1 s0 = 1 0 --> y= i2
#50 i0=0;i1=1;i2=0;i3=0;
#50 i0=0;i1=0;i2=1;i3=0;
#50 i0=0;i1=0;i2=0;i3=1;

#50 s0=1;i0=1;i1=0;i2=0;i3=0;               //s1 s0 = 1 1 --> y= i3
#50 i0=0;i1=1;i2=0;i3=0;
#50 i0=0;i1=0;i2=1;i3=0;
#50 i0=0;i1=0;i2=0;i3=1;
#50 $finish;
end
endmodule
