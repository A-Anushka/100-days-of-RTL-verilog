module nor_ga(output y,input a,input b);
nor(y,a,b);
endmodule
